`include "common/pfme_sec0.sv"
`include "common/pfme_sec1.sv"
`include "common/pfme_sec2.sv"
