../pfme_cfg_in.sv // pfme_cfg 
../pfme_a_in.sv // pfme_a 
