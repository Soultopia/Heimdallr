`include "common/pfme_cfg_in_pfme_sec0.sv"
`include "common/pfme_cfg_in_pfme_sec1.sv"
`include "common/pfme_cfg_in_pfme_sec2.sv"
