module top_test(
    input a,
    output b
);






endmodule
